module tb;
  initial begin
    $error("Hello World");
    $finish;
  end
endmodule
